���      �sklearn.linear_model._base��LinearRegression���)��}�(�fit_intercept���	normalize��
deprecated��copy_X���n_jobs�N�positive���n_features_in_�K�coef_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KKK��h�dtype����f8�����R�(K�<�NNNJ����J����K t�b�C��+?�}��t�b�	_residues�hhK ��h��R�(KK��h�C�D��m�A�t�b�rank_�K�	singular_�hhK ��h��R�(KK��h�C`��XT@�t�b�
intercept_�hhK ��h��R�(KK��h�CjԲ>�Q-A�t�b�_sklearn_version��1.0.1�ub.