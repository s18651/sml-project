��C+     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.1�ub�n_estimators�K�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hG        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK"��h+�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C�=  �  �  �  �      �  �      N  (  6  Y  �  �  �  4  ?  �  �  a  e  z  �  �  )#  �'  q+  �+  �+  9,  �-  �t�b�
n_classes_�K"�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��h4�f8�����R�(Kh8NNNJ����J����K t�b�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<h(�scalar���h4�i8�����R�(Kh8NNNJ����J����K t�bC"       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hK�
node_count�K-�nodes�h*h-K ��h/��R�(KK-��h4�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hmhPK ��hnhPK��hohPK��hphHK��hqhHK ��hrhPK(��hshHK0��uK8KKt�b�B�	                             ڞ@�W��H�?             A@                           О@���Q��?             @������������������������       �                      @������������������������       �                     @                           �@����"�?             =@                           ��@      �?              @       
                    �@
ףp=
�?             @       	                    �@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �@gG-B���?             5@                           �@VUUUUU�?             @                           �@VUUUUU�?             @������������������������       �                     �?                           
�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           *�@�6�i�?             .@                           �@�q�q�?             @������������������������       �                     �?������������������������       �                      @       *                    j�@�q�q�?
             (@       )                    ^�@������?             "@                           6�@ܶm۶m�?             @������������������������       �                     �?                            @�@�������?             @������������������������       �                     �?!       "                    F�@�������?             @������������������������       �                     �?#       $                    J�@      �?             @������������������������       �                     �?%       &                    N�@VUUUUU�?             @������������������������       �                     �?'       (                    R�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @+       ,                    n�@�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�b�values�h*h-K ��h/��R�(KK-KK"��hH�B�/         @      �?                      @      �?      �?      @      @       @              �?       @              �?      �?      �?      �?      �?      �?      �?      �?      �?                      �?                               @               @      �?               @                                                      @                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                              �?                      @      �?      �?              @       @              �?       @              �?      �?      �?      �?      �?      �?      �?      �?      �?                      �?                               @               @      �?                      �?                                                      @       @                                                      �?                              �?                                                                                                                      �?                                                               @                                                      �?                              �?                                                                                                                      �?                                                               @                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                      �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                              @                                                                                                                                                                                                                                              @      �?      �?                                      �?       @              �?      �?              �?      �?      �?              �?      �?                      �?                               @               @      �?                                              @      �?      �?                                                                                      �?                                                                                                                                                                              �?      �?                                                                                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                      �?                                                                                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                      �?       @              �?      �?                      �?      �?              �?      �?                      �?                               @               @      �?                                                                                                      �?       @                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                              �?      �?                      �?      �?              �?      �?                      �?                               @               @      �?                                                                                                                              �?      �?                      �?      �?              �?      �?                      �?                               @                                                                                                                                                      �?      �?                      �?      �?              �?      �?                      �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                      �?      �?                      �?      �?                      �?                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                      �?                      �?      �?                      �?                      �?                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                      �?                      �?      �?                                              �?                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?                      �?                                                      �?                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                      �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                               @      �?                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK/hdh*h-K ��h/��R�(KK/��hk�BH
         ,                    b�@�8�G�V�?             A@       )                    R�@��8��8�?             >@                           Ԟ@	j*D�?             :@������������������������       �                      @                           �@      �?             8@                           ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @	                           ��@p��&%��?             5@
                           �@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �@?,R�n�?             2@                           ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �@�6�i�?             .@                           �@VUUUUU�?             @                           �@VUUUUU�?             @������������������������       �                     �?                           
�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �@�q�q�?	             "@������������������������       �                     �?                           �@      �?              @������������������������       �                     �?                           $�@ܶm۶m�?             @������������������������       �                     �?                            ,�@�������?             @������������������������       �                     �?!       "                    6�@�������?             @������������������������       �                     �?#       $                    @�@      �?             @������������������������       �                     �?%       &                    F�@VUUUUU�?             @������������������������       �                     �?'       (                    L�@      �?              @������������������������       �                     �?������������������������       �                     �?*       +                    Z�@      �?             @������������������������       �                     @������������������������       �                     �?-       .                    h�@      �?             @������������������������       �                     @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK/KK"��hH�B�1         @                      �?              �?      �?               @      �?       @      @              �?      �?              �?      �?      �?      �?              �?      �?      �?       @      @              �?      �?              @      �?              �?       @                      �?              �?      �?               @      �?       @      @              �?      �?              �?      �?      �?      �?              �?      �?      �?       @      @              �?      �?                                      �?       @                      �?              �?      �?               @      �?       @      @              �?      �?              �?      �?      �?      �?              �?      �?      �?       @                      �?      �?                                               @                                                                                                                                                                                                                                                                                                      �?              �?      �?               @      �?       @      @              �?      �?              �?      �?      �?      �?              �?      �?      �?       @                      �?      �?                                                                      �?                                                       @                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                      �?      �?               @      �?              @              �?      �?              �?      �?      �?      �?              �?      �?      �?       @                      �?      �?                                                                                                                      �?                                                                                                                       @                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                      �?      �?               @                      @              �?      �?              �?      �?      �?      �?              �?      �?      �?                              �?      �?                                                                                                               @                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                               @                                                                                                                                                                                                                                                      �?      �?                                      @              �?      �?                      �?      �?      �?              �?      �?      �?                              �?      �?                                                                                      �?      �?                                      @                                              �?                                                                                                                                                                              �?      �?                                                                                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                      �?                                                                                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                              �?      �?                              �?      �?              �?      �?      �?                              �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                              �?      �?                              �?      �?              �?      �?      �?                                      �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                                      �?                              �?      �?              �?      �?      �?                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                              �?                              �?      �?              �?      �?      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                      �?                              �?      �?              �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                      �?                              �?      �?                      �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                              �?      �?                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      @                                                              �?                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                      @      �?                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                      �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK'hdh*h-K ��h/��R�(KK'��hk�B�         &                    j�@0��>���?             A@       %                    b�@-���?             ?@                            J�@n۶m۶�?             <@                           ̞@�����|�?             6@������������������������       �                      @                           Ҟ@H�z�G�?             4@������������������������       �                      @                           F�@��^B{	�?             2@	                           
�@     ��?             0@
                           �@      �?              @                           ��@9��8���?             @                           ޞ@      �?             @������������������������       �                     �?                           �@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           �@      �?              @������������������������       �                     @                           �@�������?             @������������������������       �                     �?                           ,�@      �?             @������������������������       �                     �?                           6�@VUUUUU�?             @������������������������       �                     �?                           @�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @!       "                    N�@      �?             @������������������������       �                     @#       $                    X�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK'KK"��hH�Bp)                         @                       @              �?       @      �?              �?                      �?      @              @      �?       @      �?      �?      �?      �?      �?               @                              @              @      �?                       @                       @              �?       @      �?              �?                      �?      @              @      �?       @      �?      �?      �?      �?      �?               @                              @                      �?                       @                       @              �?       @      �?              �?                      �?      @              @      �?       @      �?      �?      �?      �?      �?               @                                                      �?                       @                       @              �?       @      �?              �?                      �?                      @               @      �?      �?      �?      �?      �?               @                                                                                                                                                                                                                                                                               @                                                                               @                       @              �?       @      �?              �?                      �?                      @               @      �?      �?      �?      �?      �?                                                                                               @                                                                                                                                                                                                                                                                                                       @              �?       @      �?              �?                      �?                      @               @      �?      �?      �?      �?      �?                                                                                                                       @              �?       @      �?              �?                      �?                      @                      �?      �?      �?      �?      �?                                                                                                                       @              �?       @      �?                                                                                      �?                              �?                                                                                                                                      �?       @      �?                                                                                      �?                              �?                                                                                                                                      �?              �?                                                                                      �?                              �?                                                                                                                                      �?                                                                                                                                                                                                                                                                                              �?                                                                                      �?                              �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                      �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                               @                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                              �?                      �?                      @                              �?      �?      �?                                                                                                                                                                                                                              @                                                                                                                                                                                                                              �?                      �?                                                      �?      �?      �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                      �?      �?      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                      �?                                                      �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                      �?                                                              �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                              @                      �?                                                                                                                      �?                                                                                                                              @                                                                                                                                                                                                                                                                                                      �?                                                                                                                      �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK+hdh*h-K ��h/��R�(KK+��hk�Bh	                             Ҟ@�W��H�?             A@                           Ξ@:/����?             @                           ʞ@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @       *                    n�@�5?,R�?             ;@                           �@�<,Ԛ��?             9@	                           �@���#���?             &@
                           �@      �?              @                           ڞ@      �?             @������������������������       �                     �?                           �@VUUUUU�?             @������������������������       �                     �?                           ��@      �?              @������������������������       �                     �?������������������������       �                     �?                           
�@      �?             @������������������������       �                      @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �@�Cc}h�?
             ,@������������������������       �                      @                           ,�@      �?	             (@                           $�@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           6�@~X�<��?             "@������������������������       �                      @        !                    @�@����X�?             @������������������������       �                      @"       #                    J�@�������?             @������������������������       �                     �?$       %                    X�@      �?             @������������������������       �                     �?&       '                    d�@VUUUUU�?             @������������������������       �                     �?(       )                    j�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�t�bh�h*h-K ��h/��R�(KK+KK"��hH�B�-         @      �?      @              �?               @      �?      �?                      �?               @       @                              �?              �?       @      �?       @                       @      @      �?      �?              �?       @      �?       @              @                                                                                                                                                                                               @                                                               @                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                               @                                                               @                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                      �?                      �?               @      �?      �?                      �?               @       @                              �?              �?       @      �?       @                              @      �?      �?              �?       @      �?              �?                      �?               @      �?      �?                      �?               @       @                              �?              �?       @      �?       @                              @      �?      �?              �?              �?              �?                      �?               @      �?      �?                      �?                                                                      �?                                                      @                                                              �?                      �?               @      �?      �?                      �?                                                                      �?                                                                                                                      �?                                              �?      �?                                                                                              �?                                                                                                                                                                      �?                                                                                                                                                                                                                              �?                                                      �?                                                                                              �?                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?               @                                      �?                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                              �?                                                      �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                              @                                                                                                                                                               @       @                              �?                       @      �?       @                                      �?      �?              �?              �?                                                                                                               @                                                                                                                                                                                                                                                                                       @                              �?                       @      �?       @                                      �?      �?              �?              �?                                                                                                                                                                                               @                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                       @                                                                                                                                                                                                       @                              �?                       @      �?                                                      �?              �?              �?                                                                                                                                                                               @                                                                                                                                                                                                                       @                              �?                              �?                                                      �?              �?              �?                                                                                                                       @                                                                                                                                                                                                                                                                                                              �?                              �?                                                      �?              �?              �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                              �?                                                                                      �?              �?              �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                      �?              �?              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hK
hcK/hdh*h-K ��h/��R�(KK/��hk�BH
         
                    �@V�(��d�?             A@       	                    �@      �?              @                           ؞@
ףp=
�?             @                           ʞ@VUUUUU�?             @������������������������       �                     �?                           Ξ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @       &                    X�@XV��?             :@       %                    J�@?,R�n�?             2@                           �@     @�?             0@                           ��@{�G�z�?             @                           ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           "�@3(&ޏ�?
             &@                           �@�������?             @������������������������       �                     �?                           �@�������?             @������������������������       �                     �?                           �@      �?             @������������������������       �                     �?                           �@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?                            *�@
ףp=
�?             @������������������������       �                      @!       "                    6�@VUUUUU�?             @������������������������       �                     �?#       $                    @�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @'       (                    b�@      �?              @������������������������       �                     @)       ,                    j�@
ףp=
�?             @*       +                    f�@      �?              @������������������������       �                     �?������������������������       �                     �?-       .                    n�@�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK/KK"��hH�B�1        �?       @      �?              �?      �?      �?               @      @              �?       @              �?               @               @                      �?      �?              �?              �?      �?      �?      �?      �?       @      �?      @      �?       @      �?                                                      @                                                                                                                                      �?                                                              �?       @      �?                                                                                                                                                                                              �?                                                              �?              �?                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                              �?              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                      �?      �?      �?               @                      �?       @              �?               @               @                      �?      �?              �?                      �?      �?      �?      �?       @      �?      @                                      �?      �?      �?               @                      �?       @              �?               @               @                      �?      �?              �?                      �?      �?                                                                              �?      �?      �?               @                      �?       @              �?               @                                      �?      �?              �?                      �?      �?                                                                                                               @                                                               @                                                              �?                                                                                                                                                                                                               @                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                               @                                                                                                                                                                                                               @                                                                                                                                                                                                                                              �?      �?      �?                                      �?       @              �?                                                      �?      �?                                      �?      �?                                                                              �?      �?      �?                                      �?                                                                                                                              �?      �?                                                                                              �?                                                                                                                                                                                                                                                              �?      �?                                              �?                                                                                                                              �?      �?                                                                                      �?                                                                                                                                                                                                                                                                      �?                                                      �?                                                                                                                              �?      �?                                                                              �?                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                              �?      �?                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                              �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                               @              �?                                                      �?      �?                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                              �?                                                      �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                      �?                                                              �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                      �?      �?       @      �?      @                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                              �?      �?       @      �?                                                                                                                                                                                                                                                      �?      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                               @      �?                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                      �?        �t�bub��     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hK	hcK)hdh*h-K ��h/��R�(KK)��hk�B�         $                    R�@y�����?             A@       #                    N�@��}*_��?             ;@                           �@V-��?             9@                           �@      �?              @                           ؞@
ףp=
�?             @                           Ξ@      �?              @������������������������       �                     �?������������������������       �                     �?	       
                    ޞ@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                            �@�~Q$���?             1@                           �@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �@/����?
             ,@                           �@������?             @                           
�@      �?             @������������������������       �                     �?                           �@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           "�@4և����?             @������������������������       �                      @                            6�@
ףp=
�?             @                           &�@      �?              @������������������������       �                     �?������������������������       �                     �?!       "                    H�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @%       &                    \�@�$I�$I�?             @������������������������       �                     @'       (                    h�@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�bh�h*h-K ��h/��R�(KK)KK"��hH�B�+                �?               @      �?      �?              �?                      @      �?      �?                      �?              �?       @               @               @      �?      �?      @      �?      @       @              �?       @                              �?               @      �?      �?              �?                      @      �?      �?                      �?              �?       @               @               @      �?      �?              �?      @       @                                                      �?               @      �?      �?              �?                      @      �?      �?                      �?              �?                       @               @      �?      �?              �?      @       @                                                      �?               @                              �?                      @                                                                                                                              �?                                                                      �?               @                              �?                                                                                                                                                      �?                                                                                                                      �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                      �?                                                                                                                                                                                                                              �?               @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                              �?      �?                                              �?      �?                      �?              �?                       @               @      �?      �?                      @       @                                                                                                                                                                                                               @                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                               @                                                                                                                                              �?      �?                                              �?      �?                      �?              �?                                       @      �?                              @       @                                                                              �?      �?                                              �?                                              �?                                                                              @                                                                                      �?      �?                                              �?                                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                      �?                                                      �?                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                      �?                                                      �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                              @                                                                                                                                                      �?                      �?                                                       @      �?                                       @                                                                                                                                                                                                                                                                               @                                                                                                                                              �?                      �?                                                       @      �?                                                                                                                                                                                      �?                                                                                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                              �?                                                       @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                      @                                      �?       @                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                      �?       @                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                       @                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK)hdh*h-K ��h/��R�(KK)��hk�B�                             ��@y�����?             A@                           �@r�q��?             (@                           Ҟ@      �?              @                           Ξ@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           ؞@
ףp=
�?             @������������������������       �                      @	       
                    ޞ@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �@P*L�9�?             6@                           �@���Q��?             @������������������������       �                      @������������������������       �                     @                           �@�~Q$���?             1@                           �@{�G�z�?             @                           
�@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                            L�@�8��8��?	             (@                           *�@
ףp=
�?             @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?                           <�@�q�q�?             @������������������������       �                      @������������������������       �                     �?!       "                    Z�@������?             @������������������������       �                     @#       $                    f�@      �?             @������������������������       �                     �?%       &                    j�@VUUUUU�?             @������������������������       �                     �?'       (                    n�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK)KK"��hH�B�+        �?      �?       @      �?              �?      @       @       @      �?               @      �?                                       @      @      �?               @                      @                      �?              �?      �?      �?      �?              �?      �?       @      �?                               @              �?                                                                                                                      @                                                                              �?      �?       @      �?                               @              �?                                                                                                                                                                                                      �?               @                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                      �?              �?                               @              �?                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                              �?              �?                                              �?                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                              �?                                                              �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                      @                                                                                                                      �?      @               @                       @      �?                                       @      @      �?               @                                              �?              �?      �?      �?      �?                                                              @               @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                      �?                                               @      �?                                       @      @      �?               @                                              �?              �?      �?      �?      �?                                                      �?                                               @                                               @                                                                                                                                                                              �?                                                                                               @                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                      �?                                              @      �?               @                                              �?              �?      �?      �?      �?                                                                                                              �?                                                      �?               @                                              �?                                                                                                                                                      �?                                                                                                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?               @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                      @                                                                                      �?      �?      �?      �?                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                                      �?      �?      �?      �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                      �?              �?      �?                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                              �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hK	hcK+hdh*h-K ��h/��R�(KK+��hk�Bh	         *                    n�@ä�hJ,�?             A@                           6�@dG�+�?             ?@                           ʞ@�������?             4@������������������������       �                      @                           ؞@?,R�n�?             2@                           О@�q�q�?             @������������������������       �                     �?������������������������       �                      @	                           �@�6�i�?             .@
                           ��@      �?              @                           ޞ@      �?             @������������������������       �                     �?                           �@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?                           ��@      �?             @������������������������       �                      @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?                           �@4և����?             @������������������������       �                      @                           �@
ףp=
�?             @������������������������       �                      @                           �@VUUUUU�?             @������������������������       �                     �?                           &�@      �?              @������������������������       �                     �?������������������������       �                     �?        !                    D�@�zv��?             &@������������������������       �                     @"       %                    Z�@4և����?             @#       $                    P�@�q�q�?             @������������������������       �                     �?������������������������       �                      @&       '                    b�@      �?             @������������������������       �                      @(       )                    h�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK+KK"��hH�B�-        �?      �?              �?       @      �?               @      �?                       @              �?      @      �?       @                              �?      �?                      �?       @       @      �?                      �?      �?      @       @      �?      �?              �?       @      �?               @      �?                       @              �?      @      �?       @                              �?      �?                      �?       @       @      �?                      �?      �?               @      �?      �?              �?       @      �?               @      �?                       @              �?                       @                              �?      �?                      �?               @      �?                                                                                                                                                                                                                                                                       @                                                              �?      �?              �?       @      �?               @      �?                       @              �?                       @                              �?      �?                      �?                      �?                                                      �?                                                       @                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                              �?              �?       @      �?                      �?                       @              �?                       @                              �?      �?                      �?                      �?                                                              �?              �?              �?                      �?                                                               @                              �?                              �?                                                                                      �?              �?                                                                                                                                      �?                              �?                                                                                                      �?                                                                                                                                                                                                                                                              �?                                                                                                                                                      �?                              �?                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                                      �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                      �?                      �?                                                               @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                      �?                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                       @                                                       @              �?                                                              �?                                              �?                                                                                       @                                                                                                                                                                                                                                                                                                                                       @              �?                                                              �?                                              �?                                                                                                                                               @                                                                                                                                                                                                                                                                                              �?                                                              �?                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                              �?                                                              �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                      @      �?                                                                               @                                      �?      �?               @                                                                                                                      @                                                                                                                                                                                                                                                                                      �?                                                                               @                                      �?      �?               @                                                                                                                              �?                                                                               @                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                      �?      �?               @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                      �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK+hdh*h-K ��h/��R�(KK+��hk�Bh	         
                    ޞ@�?             A@       	                    ؞@      �?              @                           ʞ@      �?             @������������������������       �                     �?                           Ξ@VUUUUU�?             @������������������������       �                     �?                           Ҟ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                            ,�@>�Q��?             :@                           �@     ��?             0@                           ��@~X�<��?             "@                           ��@
ףp=
�?             @                           �@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �@      �?             @������������������������       �                      @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?                           �@����>4�?             @������������������������       �                     @                           �@      �?             @������������������������       �                     �?                           $�@�q�q�?             @������������������������       �                      @������������������������       �                     �?!       "                    6�@�������?             $@������������������������       �                     @#       (                    X�@4և����?             @$       '                    L�@      �?             @%       &                    B�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @)       *                    d�@�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK+KK"��hH�B�-        �?      �?      �?      @              �?              �?       @              �?      �?              �?      �?               @               @      �?              @              �?      �?              �?      @       @      �?                               @      �?              �?      @                              �?                                                                                                                                                      �?                                                              �?              �?                                      �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                              �?                                                              �?              �?                                      �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                              �?                                      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                              �?                              �?                       @              �?      �?              �?      �?               @               @      �?              @              �?      �?                      @       @      �?                               @              �?                              �?                       @              �?      �?              �?                       @                                                      �?      �?                      @       @                                                      �?                              �?                       @              �?      �?                                       @                                                              �?                                                                                      �?                                                                      �?                                               @                                                              �?                                                                                      �?                                                                      �?                                                                                                              �?                                                                                      �?                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                              �?                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                               @                                                                                                                                                                                      �?                       @                      �?                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                      �?                                              �?                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                              �?                                                                              �?                              @       @                                                                                                                                                                                                                                                                      @                                                                                                                                                              �?                                                                              �?                                       @                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                              �?                                       @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                      �?                                                                                                                                                                                                      �?                               @      �?              @                                                              �?                               @                                                                                                                                                                              @                                                                                                                                                                                                                      �?                               @      �?                                                                              �?                               @                                                                                                                      �?                               @      �?                                                                                                                                                                                                                                      �?                                      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                                      �?                               @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                              �?                                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK%hdh*h-K ��h/��R�(KK%��hk�B         "                    b�@0��>���?             A@                           @�@d��0u��?             >@                           Ξ@�"e����?             2@������������������������       �                      @                           Ҟ@     ��?
             0@������������������������       �                      @                           ؞@/����?	             ,@������������������������       �                      @	       
                    ��@�8��8��?             (@������������������������       �                      @                           ��@�z�G��?             $@������������������������       �                      @                           �@      �?              @������������������������       �                      @                           2�@9��8���?             @                           �@      �?             @������������������������       �                     �?                           "�@VUUUUU�?             @������������������������       �                     �?                           &�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           F�@9��8���?             (@������������������������       �                     @                           N�@      �?              @                           J�@      �?             @������������������������       �                     �?������������������������       �                     @                           R�@      �?             @������������������������       �                     �?        !                    Z�@�q�q�?             @������������������������       �                      @������������������������       �                     �?#       $                    h�@      �?             @������������������������       �                     @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK%KK"��hH�BP'         @               @       @                       @       @                       @              �?               @      @                      �?      �?                      @      �?               @              �?      �?              @      �?              �?       @               @       @                       @       @                       @              �?               @      @                      �?      �?                      @      �?               @              �?      �?                                      �?       @               @       @                       @       @                       @              �?               @                                                                      �?                              �?      �?                                               @                                                                                                                                                                                                                                                                                               @       @                       @       @                       @              �?               @                                                                      �?                              �?      �?                                                               @                                                                                                                                                                                                                                                                                       @                       @       @                       @              �?               @                                                                      �?                              �?      �?                                                                                                       @                                                                                                                                                                                                                                               @                       @                               @              �?               @                                                                      �?                              �?      �?                                                                       @                                                                                                                                                                                                                                                                                                       @                               @              �?               @                                                                      �?                              �?      �?                                                                                                                               @                                                                                                                                                                                                                                               @                                              �?               @                                                                      �?                              �?      �?                                                                                               @                                                                                                                                                                                                                                                                                                                              �?               @                                                                      �?                              �?      �?                                                                                                                                              �?                                                                                      �?                              �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                      �?                                                                                      �?                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                              �?                                                                                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                      @                      �?      �?                      @                       @                                                              �?                                                                                                                                                                                      @                                                                                                                                                                                                                      @                      �?      �?                                               @                                                              �?                                                                                                                              @                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                      �?                                                       @                                                              �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                       @                                                              �?                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                      @      �?                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                      �?                �t�bub�x     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJQY%hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK)hdh*h-K ��h/��R�(KK)��hk�B�                             Ҟ@y�����?             A@                           Ξ@z�G�z�?             @������������������������       �                     �?������������������������       �                     @                           ,�@o8���?             =@                           $�@�~Q$���?             1@                           �@/�����?             ,@                           �@N�zv�?	             &@	                           �@������?             "@
                           ڞ@ܶm۶m�?             @������������������������       �                     �?                           �@�������?             @������������������������       �                     �?                           �@�������?             @������������������������       �                     �?                           ��@      �?             @������������������������       �                     �?                           �@VUUUUU�?             @������������������������       �                     �?                           
�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           �@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                           <�@�������?             (@������������������������       �                     @                            J�@0�����?             "@������������������������       �                      @!       "                    N�@4և����?             @������������������������       �                      @#       &                    Z�@
ףp=
�?             @$       %                    R�@      �?              @������������������������       �                     �?������������������������       �                     �?'       (                    f�@�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK)KK"��hH�B�+        �?      �?      @               @      �?      �?      �?              �?      �?       @               @               @              �?      �?       @              @              @              �?                      �?                      �?               @      �?              @                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                      �?                       @      �?      �?      �?              �?      �?       @               @               @              �?      �?       @              @              @              �?                      �?                      �?               @              �?                       @      �?      �?      �?              �?      �?       @               @                              �?                                              @                                      �?                                                      �?                       @      �?      �?      �?              �?      �?       @               @                              �?                                                                                      �?                                                      �?                       @      �?      �?      �?              �?      �?       @                                              �?                                                                                                                                              �?                       @      �?      �?      �?              �?      �?                                                      �?                                                                                                                                              �?                              �?      �?      �?              �?      �?                                                      �?                                                                                                                                                                                              �?                                                                                                                                                                                                                              �?                              �?      �?                      �?      �?                                                      �?                                                                                                                                              �?                                                                                                                                                                                                                                                                                                              �?      �?                      �?      �?                                                      �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                      �?      �?                      �?                                                              �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?      �?                                                                                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                      �?                                                                                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                               @                                                                                                                      �?                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                      @                                                                                                                                                                                                               @                      �?       @              @                              �?                                              �?               @                                                                                                                                                                              @                                                                                                                                                                                                                               @                      �?       @                                              �?                                              �?               @                                                                                                                                                               @                                                                                                                                                                                                                                               @                      �?                                                      �?                                              �?               @                                                                                                                               @                                                                                                                                                                                                                                                                                                      �?                                                      �?                                              �?               @                                                                                                                                                      �?                                                      �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                              �?               @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                              �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��fbhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK+hdh*h-K ��h/��R�(KK+��hk�Bh	         $                    R�@h+�v:�?             A@                           2�@�<,Ԛ��?             9@       
                    �@q=
ףp�?             4@       	                    �@�q�q�?             @                           ��@      �?             @                           Ҟ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           
�@�Cc}h�?             ,@                           �@������?             @                           ��@      �?             @������������������������       �                     �?                           ��@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �@����X�?             @                           �@      �?             @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           "�@VUUUUU�?             @������������������������       �                     �?                           &�@      �?              @������������������������       �                     �?������������������������       �                     �?        !                    @�@{�G�z�?             @������������������������       �                      @"       #                    J�@�q�q�?             @������������������������       �                      @������������������������       �                     �?%       &                    Z�@��"e���?             "@������������������������       �                     @'       (                    d�@�8��8��?             @������������������������       �                     @)       *                    l�@�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK+KK"��hH�B�-                                �?              @      �?              �?               @      �?      �?       @       @              �?      �?      �?              �?               @      �?       @      @      �?              �?       @                      �?      @                              �?              @      �?              �?               @      �?      �?       @       @              �?      �?      �?              �?               @      �?       @              �?              �?                                                                      �?              @      �?              �?               @      �?      �?       @                      �?      �?                      �?                      �?       @              �?              �?                                                                      �?                                                       @                                                                                                               @              �?                                                                                      �?                                                       @                                                                                                                              �?                                                                                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                              �?                                                                                      �?                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                      @      �?              �?                      �?      �?       @                      �?      �?                      �?                      �?                                      �?                                                                                      @      �?              �?                                                              �?                              �?                                                                                                                                                              �?              �?                                                              �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                              �?              �?                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                              �?              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                              �?      �?       @                              �?                                              �?                                      �?                                                                                                                                      �?               @                              �?                                                                                                                                                                                                                              �?                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                      �?                                                                                      �?                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                              �?                                                                                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                       @                              �?                               @                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                              �?                               @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                      @                               @                      �?      @                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                               @                      �?      @                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                               @                      �?                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ$�phG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK)hdh*h-K ��h/��R�(KK)��hk�B�                             ؞@�M���?             A@������������������������       �                     @                           
�@��^����?             ?@                           �@
ףp=
�?             $@       
                    �@VUUUUU�?             @                           �@VUUUUU�?             @������������������������       �                     �?       	                    ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @                           �@^�u]�u�?             5@                           �@�q�q�?             @                           �@      �?             @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           R�@�q�q�?             .@                           N�@������?             @                           2�@      �?             @������������������������       �                     �?                           F�@VUUUUU�?             @������������������������       �                     �?                           J�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       "                    b�@      �?              @        !                    Z�@�q�q�?             @������������������������       �                     �?������������������������       �                      @#       &                    j�@
ףp=
�?             @$       %                    f�@�q�q�?             @������������������������       �                     �?������������������������       �                      @'       (                    n�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK)KK"��hH�B�+                                        �?      @      @              �?      �?                               @              �?              �?      @      �?                      �?              �?      �?      @       @      �?       @      �?      �?      �?       @                                                                                                                                                                                                                      @                                                                                              �?      @      @              �?      �?                               @              �?              �?      @      �?                      �?              �?      �?               @      �?       @      �?      �?      �?       @                                              @      @              �?      �?                                                                                                                      �?                                                                                                                              @              �?      �?                                                                                                                      �?                                                                                                                                              �?      �?                                                                                                                      �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                      �?                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                              �?                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                      �?                                                                       @              �?              �?      @      �?                      �?                      �?               @      �?       @      �?      �?      �?       @                                      �?                                                                       @                              �?                                                                               @                                                                                      �?                                                                                                      �?                                                                               @                                                                                      �?                                                                                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                               @                                                                                                                                                                                                                                                                                              �?                      @      �?                      �?                      �?                      �?       @      �?      �?      �?       @                                                                                                                              �?                      @      �?                      �?                                              �?                                                                                                                                                                      �?                              �?                      �?                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                      �?                              �?                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                      �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                      �?                               @      �?      �?      �?       @                                                                                                                                                                                                              �?                                                               @                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                               @      �?      �?      �?                                                                                                                                                                                                                                                       @      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                              �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJW:+LhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hK
hcK'hdh*h-K ��h/��R�(KK'��hk�B�                             ��@�|�l��?             A@                           ؞@h/�����?             "@                           Ξ@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @                           �@\ A�c��?             9@������������������������       �                      @	                            N�@��Ҍ��?             7@
                           �@?��M��?             1@                           �@{�G�z�?             @                           ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           
�@      �?	             (@������������������������       �                      @                           �@��Q���?             $@                           �@      �?             @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �@9��8���?             @������������������������       �                      @                           *�@      �?             @������������������������       �                     �?                           :�@VUUUUU�?             @������������������������       �                     �?                           H�@      �?              @������������������������       �                     �?������������������������       �                     �?!       "                    R�@VUUUUU�?             @������������������������       �                     @#       $                    Z�@VUUUUU�?             @������������������������       �                     �?%       &                    b�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK'KK"��hH�Bp)                                @      �?       @       @       @       @               @       @      �?                      �?      �?      �?      @                      �?      �?                      �?       @       @                      �?                      �?                              @                               @                                                                                                                                                       @                                                                                                                       @                                                                                                                                                       @                                                                                                                                                                                                                                                                               @                                                                                                                       @                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                      �?       @       @               @               @       @      �?                      �?      �?      �?      @                      �?      �?                      �?               @                      �?                      �?                                                                                       @                                                                                                                                                                                                                              �?       @       @               @                       @      �?                      �?      �?      �?      @                      �?      �?                      �?               @                      �?                      �?                                      �?       @       @               @                       @      �?                      �?      �?      �?                              �?      �?                                       @                                                                                                       @               @                                                              �?                                                                                                                                                                                                               @                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                               @                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                              �?       @                                               @      �?                      �?              �?                              �?      �?                                       @                                                                                               @                                                                                                                                                                                                                                                                      �?                                                       @      �?                      �?              �?                              �?      �?                                       @                                                                                      �?                                                       @                                              �?                                                                                                                                                                      �?                                                                                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                      �?                      �?                                              �?      �?                                       @                                                                                                                                                                                                                                                                               @                                                                                                                                                      �?                      �?                                              �?      �?                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                              �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                              �?                                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                      @                                                      �?                                      �?                      �?                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                      �?                                      �?                      �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                      �?                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                      �?                        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJF<KdhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK%hdh*h-K ��h/��R�(KK%��hk�B         $                    j�@0��>���?             A@       #                    Z�@-���?             ?@       "                    N�@n۶m۶�?             <@       !                    J�@��j+���?             9@                           :�@�����|�?             6@                           ʞ@l~X�<�?             2@������������������������       �                      @                           "�@      �?             0@	                           �@/�����?             ,@
                           ؞@�q�q�?
             (@                           Ҟ@      �?             @                           Ξ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �@      �?              @                           ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �@�������?             @������������������������       �                     �?                           �@      �?             @������������������������       �                     �?                           ��@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                            F�@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK%KK"��hH�BP'        �?              �?      �?              �?               @              �?       @       @                              @      �?              @      �?      �?       @      @              �?               @                              @              @              �?              �?      �?              �?               @              �?       @       @                              @      �?              @      �?      �?       @      @              �?               @                              @                              �?              �?      �?              �?               @              �?       @       @                              @      �?              @      �?      �?       @      @              �?               @                                                              �?              �?      �?              �?               @              �?       @       @                              @      �?                      �?      �?       @      @              �?               @                                                              �?              �?      �?              �?               @              �?       @       @                                      �?                      �?      �?       @      @              �?               @                                                              �?              �?      �?              �?               @              �?       @       @                                      �?                              �?       @                      �?               @                                                                                                                                                                                                                                                                               @                                                              �?              �?      �?              �?               @              �?       @       @                                      �?                              �?       @                      �?                                                                              �?              �?      �?              �?               @              �?       @       @                                      �?                              �?                              �?                                                                              �?              �?      �?              �?               @              �?       @                                              �?                              �?                              �?                                                                              �?              �?                                       @                                                                                                                                                                                                                      �?              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                              �?              �?                              �?       @                                              �?                              �?                              �?                                                                                                      �?                                                       @                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                      �?                              �?                                                      �?                              �?                              �?                                                                                                                                                      �?                                                                                                                                                                                                                                              �?                                                                                      �?                              �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                      �?                                                                                      �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                      �?                                                                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                              �?                      @                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                              @        �t�bub��(     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJؽ�hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK/hdh*h-K ��h/��R�(KK/��hk�BH
         .                    Z�@�E��'s�?             A@       )                    F�@     `�?             @@       "                    $�@�����?             ;@                           Ҟ@p��&%��?             5@                           ̞@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �@?,R�n�?             2@	                           �@�6�i�?             .@
                           ��@�q�q�?
             (@                           ��@����X�?             @                           ؞@�������?             @������������������������       �                     �?                           ��@      �?             @������������������������       �                     �?                           �@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �@
ףp=
�?             @������������������������       �                      @                           �@VUUUUU�?             @������������������������       �                     �?                           
�@      �?              @������������������������       �                     �?������������������������       �                     �?                           �@�q�q�?             @������������������������       �                      @������������������������       �                     �?        !                    �@�q�q�?             @������������������������       �                      @������������������������       �                     �?#       $                    ,�@VUUUUU�?             @������������������������       �                     @%       &                    6�@VUUUUU�?             @������������������������       �                     �?'       (                    @�@      �?              @������������������������       �                     �?������������������������       �                     �?*       +                    J�@{�G�z�?             @������������������������       �                      @,       -                    P�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�t�bh�h*h-K ��h/��R�(KK/KK"��hH�B�1                         @      �?       @      �?      �?      �?       @              �?      �?               @      �?       @       @      �?               @      �?      �?      �?      @      �?      �?      �?              �?                                       @                       @      �?       @      �?      �?      �?       @              �?      �?               @      �?       @       @      �?               @      �?      �?      �?      @      �?      �?      �?              �?                                                               @      �?       @      �?      �?      �?       @              �?      �?               @      �?               @      �?                      �?      �?      �?      @      �?              �?              �?                                                               @      �?       @      �?      �?      �?       @              �?      �?               @                       @      �?                      �?                              �?              �?              �?                                                               @                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                               @                                                                                                                                                                                                                                                                                      �?       @      �?      �?      �?       @              �?      �?               @                       @      �?                      �?                              �?                              �?                                                                      �?       @      �?      �?      �?       @              �?      �?                                       @      �?                      �?                              �?                                                                                                      �?              �?      �?      �?       @              �?                                               @      �?                      �?                              �?                                                                                                      �?                              �?                      �?                                               @                              �?                              �?                                                                                                      �?                              �?                      �?                                                                              �?                              �?                                                                                                                                      �?                                                                                                                                                                                                                                              �?                                                      �?                                                                              �?                              �?                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?                                                                              �?                              �?                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                              �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                               @                                                                                                                                                                                      �?      �?               @                                                                      �?                                                                                                                                                                                                       @                                                                                                                                                                                                                                                      �?      �?                                                                                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                      �?                                                                                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                       @                                                      �?                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                               @                                                                                                                      �?                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                              �?                                                      �?      �?      @                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                      �?                                                      �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                      �?                                                              �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                       @                               @                                              �?                                                                                                                                                                                                                               @                                                                                                                                                                                                                                               @                                                                              �?                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                               @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJX��vhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK1hdh*h-K ��h/��R�(KK1��hk�B�
                             ʞ@�E��'s�?             A@������������������������       �                     @                           �@NZ��Yo�?             ?@                           �@������?             @                           Ξ@      �?             @������������������������       �                     �?                           Ҟ@VUUUUU�?             @������������������������       �                     �?	       
                    ڞ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       .                    j�@�q�q�?             8@       +                    b�@y'�L��?             5@                           �@�Kh/��?             2@                           �@      �?              @                           ��@�������?             @������������������������       �                     �?                           ��@�������?             @������������������������       �                     �?                           �@      �?             @������������������������       �                     �?                           �@VUUUUU�?             @������������������������       �                     �?                           
�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           $�@��Q���?             $@������������������������       �                      @       "                    @�@      �?              @        !                    2�@�q�q�?             @������������������������       �                     �?������������������������       �                      @#       $                    H�@�������?             @������������������������       �                     �?%       &                    N�@      �?             @������������������������       �                     �?'       (                    R�@VUUUUU�?             @������������������������       �                     �?)       *                    Z�@      �?              @������������������������       �                     �?������������������������       �                     �?,       -                    f�@�q�q�?             @������������������������       �                      @������������������������       �                     �?/       0                    n�@�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK1KK"��hH�B4        �?      �?      �?               @      �?      �?      �?      �?              @                               @      �?      �?      �?      �?                              �?      �?      �?      �?      @               @      �?       @       @      �?      �?                                                                                                                                                                                                                      @                                                              �?      �?      �?               @      �?      �?      �?      �?              @                               @      �?      �?      �?      �?                              �?      �?      �?      �?                       @      �?       @       @      �?      �?      �?      �?      �?                                      �?                      @                                                                                                                                                                                              �?      �?      �?                                      �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                      �?      �?                                      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                      �?                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                               @      �?      �?              �?                                               @      �?      �?      �?      �?                              �?      �?      �?      �?                       @      �?       @       @      �?      �?                                       @      �?      �?              �?                                               @      �?      �?      �?      �?                              �?      �?      �?      �?                       @      �?       @                      �?                                       @      �?      �?              �?                                               @      �?      �?      �?      �?                              �?      �?      �?      �?                       @                                      �?                                       @      �?      �?              �?                                                              �?      �?                                                      �?                                                                                                                      �?      �?              �?                                                              �?      �?                                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                      �?      �?              �?                                                              �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                      �?      �?              �?                                                                      �?                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                      �?      �?                                                                                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                      �?                                                                                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                               @      �?                      �?                              �?      �?              �?                       @                                      �?                                                                                                                                                                                                                                       @                                                                                                                                                               @      �?                      �?                              �?      �?              �?                                                              �?                                                                                                                       @                                                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                      �?                      �?                              �?                      �?                                                              �?                                                                                                                                                                                      �?                                                                                                                                                                                                                      �?                      �?                                                      �?                                                              �?                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                      �?                                                              �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?                                                              �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?       @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                               @      �?                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���EhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK-hdh*h-K ��h/��R�(KK-��hk�B�	         &                    b�@h+�v:�?             A@                           �@�X�� �?             9@                           �@���%�?
             *@                           �@)\���(�?	             $@       
                    ؞@
ףp=
�?             @                           ̞@VUUUUU�?             @������������������������       �                     �?       	                    Ҟ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �@�������?             @������������������������       �                     �?                           ��@      �?             @������������������������       �                     �?                           �@VUUUUU�?             @������������������������       �                     �?                           
�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �@      �?	             (@������������������������       �                      @                           "�@��Q���?             $@                           �@�q�q�?             @������������������������       �                     �?������������������������       �                      @       !                    J�@����X�?             @                            <�@      �?             @                           ,�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @"       #                    N�@VUUUUU�?             @������������������������       �                     �?$       %                    X�@      �?              @������������������������       �                     �?������������������������       �                     �?'       (                    f�@�<ݚ�?             "@������������������������       �                     @)       *                    j�@{�G�z�?             @������������������������       �                      @+       ,                    n�@�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK-KK"��hH�B�/                        �?       @      @      �?              �?      �?      �?               @               @              �?              �?      �?       @      �?      �?              �?                      �?      �?               @      @       @      �?      �?                      �?       @      @      �?              �?      �?      �?               @               @              �?              �?      �?       @      �?      �?              �?                      �?      �?                                              �?                      �?       @      @      �?              �?      �?      �?                                                              �?                      �?                                              �?                                                                              �?       @              �?              �?      �?      �?                                                              �?                      �?                                              �?                                                                              �?       @                              �?                                                                                                                                                      �?                                                                              �?                                      �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                              �?                                                                              �?                                      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                              �?                      �?      �?                                                              �?                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                              �?                      �?                                                                      �?                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                      �?                      �?                                                                      �?                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                      �?                                                                                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                       @               @              �?                      �?       @              �?              �?                              �?                                              �?                                                                                               @                                                                                                                                                                                                                                                                                               @              �?                      �?       @              �?              �?                              �?                                              �?                                                                                                               @                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                               @                                                                                                                                                                                                                                                                                              �?                      �?       @              �?              �?                                                                              �?                                                                                                                                                               @              �?              �?                                                                                                                                                                                                                                                              �?              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                              �?                      �?                                                                                                                      �?                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                      �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                               @      @       @      �?                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                       @               @      �?                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                               @      �?                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ:9)bhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hK	hcK+hdh*h-K ��h/��R�(KK+��hk�Bh	         (                    j�@ä�hJ,�?             A@       '                    \�@XϊF�?             >@                           �@x9/���?             <@                           �@��8��8�?             (@                           �@�����H�?             "@       	                    Ξ@9��8���?             @                           ʞ@�q�q�?             @������������������������       �                     �?������������������������       �                      @
                           Ҟ@VUUUUU�?             @������������������������       �                     �?                           ڞ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @                           �@     ��?             0@                           ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �@���%�?
             *@                           �@�Q����?             @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       "                    *�@      �?              @                           �@      �?             @������������������������       �                     �?                           �@VUUUUU�?             @������������������������       �                     �?        !                    "�@      �?              @������������������������       �                     �?������������������������       �                     �?#       $                    >�@      �?             @������������������������       �                      @%       &                    N�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @)       *                    n�@      �?             @������������������������       �                     @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK+KK"��hH�B�-         @      �?      �?              @              �?      �?       @      @      @      �?      �?                      �?              �?      �?              �?       @                                      �?      �?      �?       @              @      �?               @      �?      �?              @              �?      �?       @      @      @      �?      �?                      �?              �?      �?              �?       @                                      �?      �?      �?       @                                       @      �?      �?              @              �?      �?       @      @      @      �?      �?                      �?              �?      �?              �?       @                                      �?      �?      �?                                               @      �?      �?                                      �?              @      @                                                                                                                              �?                                                               @      �?      �?                                      �?                      @                                                                                                                              �?                                                               @      �?      �?                                      �?                                                                                                                                                      �?                                                               @                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                               @                                                                                                                                                                                                                                                                                      �?      �?                                      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                      �?                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                      @              �?               @                      �?      �?                      �?              �?      �?              �?       @                                              �?      �?                                                                                                               @                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                               @                                                                                                                                                                                                                                              @              �?                                      �?      �?                      �?              �?      �?                       @                                              �?      �?                                                                              @              �?                                                                                      �?                                                                                                                                                                                      �?                                                                                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                      �?      �?                      �?                      �?                       @                                              �?      �?                                                                                                                                      �?      �?                                                                                                                      �?      �?                                                                                                                                      �?                                                                                                                                                                                                                                                                                      �?                                                                                                                      �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                      �?                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                      �?                       @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                              �?                      �?                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                              @      �?                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�BHzhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK"��hH�B                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@�t�bh<hMhPC"       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C"       �t�bK��R�}�(hKhcK'hdh*h-K ��h/��R�(KK'��hk�B�                             �@Sbq����?             A@                           ��@�r
^N��?	             ,@                           ؞@4և����?             @                           Ξ@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �@      �?             @������������������������       �                      @	       
                    �@      �?              @������������������������       �                     �?������������������������       �                     �?                           
�@����>4�?             @������������������������       �                     @                           �@      �?             @������������������������       �                      @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?                           "�@333333�?             4@������������������������       �                     @                           *�@/����?
             ,@������������������������       �                     @       $                    f�@N�zv�?	             &@                           P�@      �?              @                           6�@      �?             @������������������������       �                     �?                           @�@VUUUUU�?             @������������������������       �                     �?                           H�@      �?              @������������������������       �                     �?������������������������       �                     �?        !                    Z�@      �?             @������������������������       �                      @"       #                    b�@      �?              @������������������������       �                     �?������������������������       �                     �?%       &                    j�@�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK'KK"��hH�Bp)        �?       @       @               @              @                              �?      �?      @              �?      �?                                              �?      �?              �?       @              �?      @       @      �?      �?              �?      �?       @       @               @              @                              �?      �?                                                                                                      �?                      �?                                                      �?       @       @                                                              �?                                                                                                              �?                                                                              �?               @                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                       @                                                                      �?                                                                                                              �?                                                                                       @                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                              �?                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                               @              @                                      �?                                                                                                                              �?                                                                                                      @                                                                                                                                                                                                                                                               @                                                      �?                                                                                                                              �?                                                                                       @                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                              �?                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                      @              �?      �?                                              �?      �?                       @                      @       @      �?      �?              �?                                                                                                                                                                                                                                      @                                                                                                                                              @              �?      �?                                              �?      �?                       @                               @      �?      �?              �?                                                                                                      @                                                                                                                                                                                                                                                                                              �?      �?                                              �?      �?                       @                               @      �?      �?              �?                                                                                                                      �?      �?                                              �?      �?                       @                                      �?                      �?                                                                                                                      �?      �?                                              �?      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                      �?      �?                                                      �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                      �?                                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                               @                                      �?                      �?                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                      �?                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                       @              �?                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                              �?                �t�bub�       hhubehhub.