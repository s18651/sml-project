��"     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.1�ub�n_estimators�K�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hG        �n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK&��h+�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C�=  �  �  �  �      �  �      7  N  (  6  Y  �  �  �  4  ?  L  �  �  a  e  z  �  �  f!  )#  �'  q+  �+  �+  9,  �-  �;  �t�b�
n_classes_�K&�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��h4�f8�����R�(Kh8NNNJ����J����K t�b�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<h(�scalar���h4�i8�����R�(Kh8NNNJ����J����K t�bC&       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hK�
node_count�K5�nodes�h*h-K ��h/��R�(KK5��h4�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hmhPK ��hnhPK��hohPK��hphHK��hqhHK ��hrhPK(��hshHK0��uK8KKt�b�B�                             �@�|�ʒ��?             C@                           �@�.k���?
             1@                           �@�r
^N��?	             ,@                           ��@�q�q�?             (@                           �@����X�?             @                           Ξ@�������?             @������������������������       �                     �?       	                    ؞@      �?             @������������������������       �                     �?
                           ��@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           ��@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @                           �@p��&%��?             5@������������������������       �                     @                           �@�E����?             2@������������������������       �                      @       *                    X�@     ��?             0@                           $�@�q�q�?	             "@������������������������       �                     �?                           *�@      �?              @������������������������       �                     �?                           .�@ܶm۶m�?             @������������������������       �                     �?        !                    4�@�������?             @������������������������       �                     �?"       #                    :�@�������?             @������������������������       �                     �?$       %                    B�@      �?             @������������������������       �                     �?&       '                    L�@VUUUUU�?             @������������������������       �                     �?(       )                    R�@      �?              @������������������������       �                     �?������������������������       �                     �?+       ,                    ^�@����X�?             @������������������������       �                      @-       .                    b�@�������?             @������������������������       �                     �?/       0                    f�@      �?             @������������������������       �                     �?1       2                    j�@VUUUUU�?             @������������������������       �                     �?3       4                    n�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�b�values�h*h-K ��h/��R�(KK5KK&��hH�B�>                                �?                       @      �?       @      �?      �?              @               @      �?              @              �?      �?      �?       @      �?              �?              �?      �?      �?      @      �?      �?      �?      �?      �?      �?       @                              �?                       @      �?       @      �?      �?              @                                      @                                       @                                              �?                                                                                                      �?                       @      �?       @      �?      �?                                                      @                                       @                                              �?                                                                                                      �?                              �?       @      �?      �?                                                      @                                       @                                              �?                                                                                                      �?                              �?              �?      �?                                                                                               @                                              �?                                                                                                      �?                              �?              �?      �?                                                                                                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                      �?                              �?              �?      �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                              �?                                              �?      �?                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                              �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                               @                                                                      @                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                               @      �?                              �?      �?      �?              �?              �?              �?              �?      @      �?      �?      �?      �?      �?      �?       @                                                                                                                                                                                                                                                      @                                                                                                                                                                               @      �?                              �?      �?      �?              �?              �?              �?              �?              �?      �?      �?      �?      �?      �?       @                                                                                                                       @                                                                                                                                                                                                                                                                                                                      �?                              �?      �?      �?              �?              �?              �?              �?              �?      �?      �?      �?      �?      �?       @                                                                                                                              �?                              �?      �?      �?              �?              �?              �?              �?              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                              �?                              �?      �?      �?              �?              �?              �?              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                              �?                              �?      �?      �?              �?                              �?              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                              �?                              �?      �?      �?              �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?                              �?      �?      �?                                              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                              �?                              �?      �?                                                      �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                              �?      �?                                                      �?                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                      �?                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                      �?      �?      �?      �?      �?       @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                      �?      �?      �?      �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?      �?      �?      �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?              �?      �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                              �?      �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                      �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hK
hcK3hdh*h-K ��h/��R�(KK3��hk�B(                             ޞ@B+K&:~�?             C@                           ؞@����>4�?             @                           Ҟ@      �?             @                           Ξ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @	       
                    �@��W64<�?             ?@������������������������       �                      @                            &�@����"�?             =@                           "�@     ��?             0@                           �@�wɃg�?
             *@                           ��@�q�q�?             @                           ��@      �?             @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           �@����X�?             @                           
�@      �?             @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @!       "                    *�@���%�?
             *@������������������������       �                     @#       .                    b�@)\���(�?	             $@$       %                    2�@�������?             @������������������������       �                     �?&       '                    @�@�������?             @������������������������       �                     �?(       )                    J�@      �?             @������������������������       �                     �?*       +                    P�@VUUUUU�?             @������������������������       �                     �?,       -                    Z�@      �?              @������������������������       �                     �?������������������������       �                     �?/       0                    f�@      �?             @������������������������       �                      @1       2                    l�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK3KK&��hH�B�<        �?       @      �?      @      �?      �?      �?       @       @      �?              �?              @      �?              �?       @       @              �?      �?                              @              �?              �?              �?      �?       @              �?      �?              �?              �?      @                               @                                                                                                                                                                                                                                                      �?              �?                                       @                                                                                                                                                                                                                                                      �?              �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                               @                      �?      �?      �?               @      �?              �?              @      �?              �?       @       @              �?      �?                              @              �?              �?              �?      �?       @              �?      �?                       @                                                                                                                                                                                                                                                                                                                                      �?      �?      �?               @      �?              �?              @      �?              �?       @       @              �?      �?                              @              �?              �?              �?      �?       @              �?      �?                                              �?      �?      �?               @      �?              �?              @      �?                       @       @                                                                                                      �?                                                                                      �?      �?      �?               @      �?              �?                      �?                       @       @                                                                                                      �?                                                                                                                       @      �?              �?                                               @                                                                                                                                                                                                                                              �?              �?                                               @                                                                                                                                                                                                                                              �?              �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                              �?      �?      �?                                                              �?                               @                                                                                                      �?                                                                                              �?      �?                                                                                               @                                                                                                                                                                                                      �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                              �?                                                                              �?                                                                                                                                      �?                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                      �?                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                      �?                              �?      �?                              @              �?              �?                      �?       @              �?      �?                                                                                                                                                                                                                      @                                                                                                                                                                                                                                      �?                              �?      �?                                              �?              �?                      �?       @              �?      �?                                                                                                                                              �?                              �?      �?                                              �?              �?                                                      �?                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                      �?                              �?      �?                                              �?                                                                      �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                      �?                              �?                                                      �?                                                                      �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                      �?                                                                      �?                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                              �?       @              �?                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                      �?                      �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hKhcK-hdh*h-K ��h/��R�(KK-��hk�B�	         $                    N�@f��.�?             C@                           :�@�������?             ;@                           �@��Q��?             4@                           �@/����?
             ,@                           �@9��8���?             @                           ʞ@      �?             @������������������������       �                     �?       	                    ֞@VUUUUU�?             @������������������������       �                     �?
                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           ��@      �?              @������������������������       �                     @                            �@
ףp=
�?             @������������������������       �                      @                           
�@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?                           &�@VUUUUU�?             @������������������������       �                     @                           *�@VUUUUU�?             @������������������������       �                     �?                           2�@      �?              @������������������������       �                     �?������������������������       �                     �?                           @�@����>4�?             @������������������������       �                     @        !                    F�@      �?             @������������������������       �                      @"       #                    J�@      �?              @������������������������       �                     �?������������������������       �                     �?%       &                    R�@*L�9��?             &@������������������������       �                     @'       ,                    h�@����>4�?             @(       +                    ^�@�Q����?             @)       *                    X�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�t�bh�h*h-K ��h/��R�(KK-KK&��hH�Bp5        �?      �?                      �?              �?                       @      �?              �?      @              @      �?       @              @      �?      �?                       @      �?      @      �?      �?      �?                                               @      @      �?      �?      �?                      �?              �?                       @      �?              �?      @              @      �?       @                      �?      �?                       @      �?      @              �?      �?                                                                      �?      �?                      �?              �?                       @      �?              �?      @                               @                              �?                              �?      @              �?      �?                                                                      �?      �?                      �?              �?                       @      �?              �?                                       @                                                                      @              �?                                                                              �?      �?                                                               @      �?                                                                                                                                              �?                                                                              �?      �?                                                                      �?                                                                                                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                              �?      �?                                                                      �?                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                      �?                                                                      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                      �?              �?                                              �?                                       @                                                                      @                                                                                                                                                                                                                                                                                                              @                                                                                                                              �?              �?                                              �?                                       @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                      �?              �?                                              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                              �?                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                      @                                                              �?                              �?                              �?                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                                              �?                              �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                              @      �?                              �?                               @                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                      �?                              �?                               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                              �?                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                      @                                                              �?                                                               @      @      �?                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                                              �?                                                               @      @      �?                                                                                                                                                                                                                              �?                                                                      @      �?                                                                                                                                                                                                                              �?                                                                              �?                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                       @                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hKhcK/hdh*h-K ��h/��R�(KK/��hk�BH
                             ʞ@(�@݈g�?             C@������������������������       �                     @       .                    j�@L�w�Z�?            �A@                           Ξ@     P�?             @@������������������������       �                      @       -                    b�@��8��8�?             >@       $                    @�@����X�?             <@       #                    :�@<��KM��?             3@	       "                    4�@e�7�
t�?             1@
                           ܞ@�*;L�?             .@                           Ҟ@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           ��@9��8���?             (@                           �@      �?             @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           ��@      �?              @������������������������       �                     �?                           
�@ܶm۶m�?             @������������������������       �                     �?                           �@�������?             @������������������������       �                     �?                           �@�������?             @������������������������       �                     �?                           "�@      �?             @������������������������       �                     �?                           *�@VUUUUU�?             @������������������������       �                     �?        !                    .�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @%       &                    F�@�2�tk~�?             "@������������������������       �                     @'       *                    P�@�q�q�?             @(       )                    J�@�q�q�?             @������������������������       �                     �?������������������������       �                      @+       ,                    X�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK/KK&��hH�B�7         @              �?                                       @      �?              �?       @      �?              �?       @       @      �?                      �?       @              �?      @      �?      �?       @      @      �?      �?               @              @                      �?                                                                                                                                                                                                                                      @                                                                               @              �?                                       @      �?              �?       @      �?              �?       @       @      �?                      �?       @              �?      @      �?      �?       @              �?      �?               @              @                      �?       @              �?                                       @      �?              �?       @      �?              �?       @       @      �?                      �?       @              �?      @      �?      �?       @              �?      �?               @                                      �?       @                                                                                                                                                                                                                                                                                                                              �?                                       @      �?              �?       @      �?              �?       @       @      �?                      �?       @              �?      @      �?      �?       @              �?      �?               @                                      �?                      �?                                       @      �?              �?       @      �?              �?       @       @      �?                      �?       @              �?      @      �?      �?       @              �?      �?                                                      �?                      �?                                       @      �?              �?       @      �?              �?       @              �?                               @              �?              �?      �?                      �?      �?                                                                              �?                                       @      �?              �?       @      �?              �?                      �?                               @              �?              �?      �?                      �?      �?                                                                              �?                                       @      �?              �?       @      �?              �?                      �?                                              �?              �?      �?                      �?      �?                                                                              �?                                       @                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                      �?              �?       @      �?              �?                      �?                                              �?              �?      �?                      �?      �?                                                                                                                                              �?       @                                                                                                                      �?                                                                                                                                                                              �?                                                                                                                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                      �?                              �?              �?                      �?                                              �?              �?                              �?      �?                                                                                                                                                                                                      �?                                                                                                                                                                                                                                      �?                              �?              �?                                                                      �?              �?                              �?      �?                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                              �?              �?                                                                      �?              �?                              �?      �?                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                              �?                                                                      �?              �?                              �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                              �?                                                                      �?              �?                              �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                      �?              �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                              �?                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                       @                              �?                              @                       @                                                                              �?                                                                                                                                                                                                      @                                                                                                                                                                                                                                               @                              �?                                                       @                                                                              �?                                                                                                                                       @                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                              �?                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                              @                        �t�bub��     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hK	hcK5hdh*h-K ��h/��R�(KK5��hk�B�                             �@\�Uo��?             C@                           
�@      �?
             0@                           �@������?	             *@                           ��@��Q���?             $@                           ��@����X�?             @                           ̞@�������?             @������������������������       �                     �?       	                    ؞@      �?             @������������������������       �                     �?
                           �@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                           "�@n,�Ra��?             6@                           �@{�G�z�?             @                           �@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @       "                    4�@e�7�
t�?             1@       !                    .�@
ףp=
�?             @                           &�@VUUUUU�?             @������������������������       �                     �?                            *�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @#       *                    N�@�q�q�?
             (@$       )                    F�@
ףp=
�?             @%       &                    :�@VUUUUU�?             @������������������������       �                     �?'       (                    @�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @+       0                    f�@����X�?             @,       /                    `�@      �?             @-       .                    X�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @1       2                    j�@VUUUUU�?             @������������������������       �                     �?3       4                    n�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK5KK&��hH�B�>                �?      �?              @              @              �?                      �?              �?       @      �?               @                       @      �?       @       @      �?      �?      �?      �?      �?      �?      �?       @      �?       @      �?      �?              �?              �?      �?              @              @              �?                      �?                                               @                                       @                              �?              �?                                                                                      �?      �?                              @              �?                      �?                                               @                                       @                              �?              �?                                                                                      �?      �?                                              �?                      �?                                               @                                       @                              �?              �?                                                                                      �?      �?                                                                      �?                                                                                       @                              �?              �?                                                                                      �?      �?                                                                      �?                                                                                                                      �?              �?                                                                                                                                                                                                                                                                                                              �?                                                                                      �?      �?                                                                      �?                                                                                                                      �?                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                                              �?                                                                                                                      �?                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                              �?                                                                       @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                                                      �?       @      �?                                       @      �?               @      �?      �?              �?              �?      �?       @      �?       @      �?      �?              �?                                                                                                                       @                                                                                                                              �?       @                                                                                                                                                                       @                                                                                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                              �?              �?                                       @      �?               @      �?      �?              �?              �?                      �?       @      �?      �?              �?                                                                                                              �?                                                                               @              �?                              �?                                                                                                                                                                              �?                                                                                              �?                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                              �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                              �?                                       @      �?                      �?                      �?                                      �?       @      �?      �?              �?                                                                                                                              �?                                       @      �?                      �?                                                                                                                                                                                                                                      �?                                              �?                      �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                              �?                                                                      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                      �?                                      �?       @      �?      �?              �?                                                                                                                                                                                                                              �?                                               @                              �?                                                                                                                                                                                                                              �?                                                                              �?                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                      �?              �?      �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                              �?      �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                      �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hK	hcK-hdh*h-K ��h/��R�(KK-��hk�B�	                             ޞ@�����?             C@                           ؞@��E���?             "@                           Ξ@      �?             @������������������������       �                     �?                           Ҟ@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @	                           ��@!��w���?             =@
                           �@      �?              @                           �@      �?             @������������������������       �                     �?                           �@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                           �@^�u]�u�?             5@                           
�@�8��8��?             @                            �@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                            �@�6�i�?             .@                           �@      �?             @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @       "                    .�@N�zv�?	             &@       !                    *�@      �?             @                            &�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @#       &                    L�@����X�?             @$       %                    <�@�q�q�?             @������������������������       �                     �?������������������������       �                      @'       (                    X�@      �?             @������������������������       �                     �?)       *                    b�@VUUUUU�?             @������������������������       �                     �?+       ,                    j�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK-KK&��hH�Bp5        �?      �?       @      @               @              �?                       @      @      �?      �?       @                              @      �?       @              �?      �?              �?      �?                       @      �?                      �?              �?      �?              �?               @      @                              �?                                                                                                                                                                                                                                                      �?               @                                      �?                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                               @                                      �?                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                              �?                               @                                       @      @      �?      �?       @                              @      �?       @              �?      �?              �?      �?                       @      �?                      �?              �?      �?                      �?                                                                       @      @                                                                                                                      �?                                                                                                      �?                                                                       @                                                                                                                              �?                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                              �?                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                      @                                                                                                                                                                                                                                                               @                                                      �?      �?       @                              @      �?       @              �?      �?              �?                               @      �?                      �?              �?      �?                                                       @                                                                                                      @                              �?                                                                                                                                                                       @                                                                                                                                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                              �?      �?       @                                      �?       @                      �?              �?                               @      �?                      �?              �?      �?                                                                                                              �?               @                                                                                                                              �?                                                                                                                                                              �?                                                                                                                                              �?                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                      �?                                              �?       @                      �?              �?                               @                              �?              �?      �?                                                                                                                      �?                                                                                              �?                               @                                                                                                                                                                              �?                                                                                              �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                              �?       @                      �?                                                                              �?              �?      �?                                                                                                                                                                               @                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                      �?                                                                                                              �?              �?      �?                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                              �?              �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                      �?              �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                              �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hK	hcK+hdh*h-K ��h/��R�(KK+��hk�Bh	                             �@f��.�?             C@                           ڞ@�q�q�?             @������������������������       �                      @������������������������       �                     @       &                    b�@     �?             @@                           F�@\ A�c��?             9@                           @�@ҳ�wY;�?             1@                           ��@�6�i�?             .@	                           ��@      �?             @
                           ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           &�@N�zv�?	             &@                           �@����X�?             @                           �@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?                           �@      �?             @������������������������       �                      @                            �@      �?              @������������������������       �                     �?������������������������       �                     �?                           ,�@      �?             @������������������������       �                      @                           6�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @        !                    N�@      �?              @������������������������       �                     @"       #                    X�@{�G�z�?             @������������������������       �                      @$       %                    ^�@�q�q�?             @������������������������       �                     �?������������������������       �                      @'       (                    f�@������?             @������������������������       �                     @)       *                    l�@      �?             @������������������������       �                     @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK+KK&��hH�B3                @                              �?      �?       @      �?                      �?       @      �?      �?      �?               @                      @              �?      �?       @       @               @                                      @      @              �?       @      �?              @                                               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                              �?      �?              �?                      �?       @      �?      �?      �?               @                      @              �?      �?       @       @               @                                      @      @              �?       @      �?                                              �?      �?              �?                      �?       @      �?      �?      �?               @                      @              �?      �?       @       @               @                                                                       @      �?                                              �?      �?              �?                      �?       @      �?      �?      �?               @                                      �?      �?       @       @                                                                                                                                              �?      �?              �?                      �?       @      �?      �?      �?               @                                      �?      �?               @                                                                                                                                                                                              �?                                               @                                      �?                                                                                                                                                                                                                      �?                                                                                      �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                              �?      �?              �?                               @      �?      �?      �?                                                              �?               @                                                                                                                                              �?      �?              �?                               @      �?      �?                                                                                                                                                                                                                                      �?      �?              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                      �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                       @      �?      �?                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                      �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                              �?                                                              �?               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                              �?                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                              @                                                       @                                                                       @      �?                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                                                       @                                                                       @      �?                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                                       @      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                              @      @              �?                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                      @                      �?                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                      �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hKhcK/hdh*h-K ��h/��R�(KK/��hk�BH
                             ؞@�5��P�?             C@                           Ξ@      �?             @������������������������       �                     �?������������������������       �                     @       $                    4�@ä�hJ,�?             A@                           ޞ@x��J��?             7@������������������������       �                      @       !                    &�@gG-B���?             5@	                           �@l~X�<�?             2@
                           �@2Tv���?             .@                           �@��Q���?             $@                           �@      �?              @                           �@      �?             @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           ��@      �?             @������������������������       �                     �?                           ��@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �@{�G�z�?             @������������������������       �                      @                           �@�q�q�?             @������������������������       �                      @������������������������       �                     �?                            "�@�q�q�?             @������������������������       �                      @������������������������       �                     �?"       #                    ,�@�q�q�?             @������������������������       �                      @������������������������       �                     �?%       &                    :�@�ˠT�?             &@������������������������       �                     @'       (                    D�@������?             @������������������������       �                     @)       *                    N�@      �?             @������������������������       �                     �?+       ,                    R�@VUUUUU�?             @������������������������       �                     �?-       .                    b�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK/KK&��hH�B�7                �?               @       @      �?              @      �?              �?      �?       @      �?      �?      @      �?      �?              �?              @              �?               @       @      �?      �?               @       @                              �?                                                                              @                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                      @                                                                                                                                                                                                                                                              �?               @       @      �?                      �?              �?      �?       @      �?      �?      @      �?      �?              �?              @              �?               @       @      �?                       @       @                              �?                              �?               @       @      �?                      �?              �?      �?       @      �?      �?                      �?                                              �?               @       @                               @       @                                                                               @                                                                                                                                                                                                                                                                                              �?                       @      �?                      �?              �?      �?       @      �?      �?                      �?                                              �?               @       @                               @       @                                                              �?                       @      �?                      �?              �?      �?       @      �?      �?                      �?                                                                       @                               @       @                                                              �?                       @      �?                      �?              �?      �?       @              �?                      �?                                                                       @                               @                                                                      �?                       @      �?                      �?              �?      �?                                              �?                                                                       @                                                                                                      �?                              �?                      �?              �?      �?                                              �?                                                                       @                                                                                                      �?                                                                      �?                                                                                                                               @                                                                                                      �?                                                                      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                      �?                      �?                      �?                                              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                              �?                      �?                                                                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                              �?                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                                               @              �?                                                                                                                               @                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                              �?                                                                                                                               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                              �?               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              @      �?                      �?              @                                              �?                                                              �?                                                                                                                                                                                              @                                                                                                                                                                                                                                                              @      �?                      �?                                                              �?                                                              �?                                                                                                                                              @                                                                                                                                                                                                                                                                                                                      �?                      �?                                                              �?                                                              �?                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?                                                              �?                                                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                �t�bub�      hhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hK
hcK/hdh*h-K ��h/��R�(KK/��hk�BH
         ,                    h�@����~E�?             C@       '                    P�@�?             A@                           ��@!��w���?             =@                           �@�T�x?r�?             &@                           ؞@9��8���?             @                           Ξ@�q�q�?             @������������������������       �                     �?������������������������       �                      @	       
                    �@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?                           ��@���Q��?             @������������������������       �                     @������������������������       �                      @                           
�@�q�q�?             2@                           �@z�G�z�?             @������������������������       �                     �?������������������������       �                     @                           �@�wɃg�?
             *@                           �@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           $�@��Q���?             $@                           �@�q�q�?             @������������������������       �                     �?������������������������       �                      @       $                    F�@����X�?             @                           ,�@      �?             @������������������������       �                     �?        !                    4�@VUUUUU�?             @������������������������       �                     �?"       #                    >�@      �?              @������������������������       �                     �?������������������������       �                     �?%       &                    J�@�q�q�?             @������������������������       �                      @������������������������       �                     �?(       )                    X�@�Q����?             @������������������������       �                     @*       +                    `�@      �?              @������������������������       �                     �?������������������������       �                     �?-       .                    n�@      �?             @������������������������       �                     @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK/KK&��hH�B�7        �?      �?       @               @      @                      �?      �?              @      �?                              �?       @      �?               @      �?              �?      �?      �?      �?      @                               @              �?      @      �?              �?      �?      �?       @               @      @                      �?      �?              @      �?                              �?       @      �?               @      �?              �?      �?      �?      �?      @                               @              �?                              �?      �?      �?       @               @      @                      �?      �?              @      �?                              �?       @      �?               @      �?              �?      �?      �?      �?                                       @                                                      �?      �?       @                                                      �?              @                                               @                                                                      �?                                                                                              �?      �?       @                                                      �?                                                                                                                                      �?                                                                                              �?               @                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                      �?                                                              �?                                                                                                                                      �?                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                      �?                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                      @                                               @                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                       @      @                      �?                              �?                              �?              �?               @      �?              �?      �?      �?                                               @                                                                                              @                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                       @                                                              �?                              �?              �?               @      �?              �?      �?      �?                                               @                                                                                       @                                                                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                              �?                              �?                               @      �?              �?      �?      �?                                               @                                                                                                                                                      �?                                                                                                                                                       @                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                      �?                               @      �?              �?      �?      �?                                                                                                                                                                                                                                                                              �?              �?      �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?              �?      �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                              �?                      �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                              �?                               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                      @                                              �?                              �?                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                              �?                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                      @      �?                                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                      �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hK	hcK)hdh*h-K ��h/��R�(KK)��hk�B�         "                    L�@f��.�?             C@                           (�@���ϭ�?             =@                            �@��Q��?             4@                           �@?��M��?             1@                           �@�Cc}h�?
             ,@                           ��@~X�<��?             "@                           �@����X�?             @                           ֞@      �?             @	       
                    Ξ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �@VUUUUU�?             @������������������������       �                     �?                           ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           
�@{�G�z�?             @������������������������       �                      @                           �@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                           2�@�<ݚ�?             "@������������������������       �                     @                           >�@{�G�z�?             @������������������������       �                      @        !                    F�@�q�q�?             @������������������������       �                      @������������������������       �                     �?#       $                    Z�@B{	�%��?             "@������������������������       �                     @%       &                    f�@VUUUUU�?             @������������������������       �                      @'       (                    j�@      �?             @������������������������       �                      @������������������������       �                      @�t�bh�h*h-K ��h/��R�(KK)KK&��hH�B�0        �?              �?       @      �?       @                       @      �?              �?       @      @      �?                               @      @      �?       @      �?               @                                      @                       @       @       @                              �?              �?       @      �?       @                       @      �?              �?       @      @      �?                               @              �?       @      �?               @                                      @                                                                      �?              �?       @      �?       @                       @      �?              �?       @      @      �?                               @                              �?                                                                                                                              �?              �?       @      �?       @                       @      �?              �?       @              �?                               @                              �?                                                                                                                              �?              �?       @      �?       @                       @      �?              �?                                                       @                              �?                                                                                                                              �?              �?       @                                       @      �?              �?                                                                                      �?                                                                                                                              �?              �?       @                                              �?              �?                                                                                      �?                                                                                                                              �?              �?       @                                                                                                                                                                                                                                                                                      �?              �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                              �?              �?                                                                                      �?                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                              �?                                                                                      �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                               @                                                                                                                                                                                                                                                                              �?       @                                                                                                       @                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                      �?                                                                                                               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                               @              �?                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                                                      �?       @                       @                                      @                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                      �?       @                       @                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                      �?                               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      @                                                                                                       @       @       @                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                                                                                                       @       @       @                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                       @               @                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                               @                        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJQY%hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hK
hcK-hdh*h-K ��h/��R�(KK-��hk�B�	                             Ξ@����~E�?             C@������������������������       �                     @                           :�@��#��2�?            �A@                           "�@l~X�<�?             2@                           �@2Tv���?             .@                           �@      �?	             (@                           �@~X�<��?             "@                           �@9��8���?             @	       
                    Ҟ@VUUUUU�?             @������������������������       �                     �?                           ؞@      �?              @������������������������       �                     �?������������������������       �                     �?                           ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           ,�@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           F�@:߄*�u�?	             1@������������������������       �                     @                            J�@�	j*D�?             *@������������������������       �                      @!       "                    N�@�T�x?r�?             &@������������������������       �                      @#       $                    R�@�����H�?             "@������������������������       �                      @%       &                    Z�@������?             @������������������������       �                     @'       (                    b�@      �?             @������������������������       �                     �?)       *                    f�@VUUUUU�?             @������������������������       �                     �?+       ,                    l�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK-KK&��hH�Bp5        @              �?      �?       @               @      �?      �?       @                      �?              �?               @              �?       @       @                      �?      @       @              @                       @              �?      �?              �?      �?              @                                                                                                                                                                                                                                                                                                                              �?      �?       @               @      �?      �?       @                      �?              �?               @              �?       @       @                      �?      @       @              @                       @              �?      �?              �?      �?                              �?      �?       @               @      �?      �?       @                      �?              �?                              �?                                      �?               @                                       @                                                                              �?      �?       @               @      �?      �?       @                      �?              �?                              �?                                                                                               @                                                                              �?      �?       @               @      �?      �?       @                      �?                                              �?                                                                                                                                                                              �?      �?                       @      �?      �?       @                                                                      �?                                                                                                                                                                              �?      �?                              �?      �?       @                                                                                                                                                                                                                                                      �?      �?                              �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                      �?                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                      �?       @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                               @                                                                                              �?                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                               @                                                              �?                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                              �?                                                                                                                               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                      �?               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                       @                       @       @                              @                      @                                      �?      �?              �?      �?                                                                                                                                                                                                              @                                                                                                                                                                                                                                               @                       @       @                                                      @                                      �?      �?              �?      �?                                                                                                                                                                               @                                                                                                                                                                                                                                                                               @                       @                                                              @                                      �?      �?              �?      �?                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                       @                                                              @                                      �?      �?              �?      �?                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                                              @                                      �?      �?              �?      �?                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                                      �?      �?              �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?      �?              �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                      �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��fbhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hK	hcK3hdh*h-K ��h/��R�(KK3��hk�B(         2                    n�@B+K&:~�?             C@                           �@A��Oru�?            �A@                           ޞ@�����H�?             "@                           ؞@������?             @                           ʞ@      �?             @������������������������       �                     �?                           Ξ@VUUUUU�?             @������������������������       �                     �?	       
                    Ҟ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @                           �@XV��?             :@                           �@>
ףp=�?             $@                           
�@����X�?             @                           �@�������?             @������������������������       �                     �?                           �@      �?             @������������������������       �                     �?                           ��@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @       #                    :�@      �?             0@       "                    2�@�q�q�?             @       !                    *�@      �?             @                            $�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @$       )                    T�@��Q���?             $@%       (                    J�@      �?             @&       '                    B�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @*       +                    ^�@9��8���?             @������������������������       �                      @,       -                    b�@      �?             @������������������������       �                     �?.       /                    f�@VUUUUU�?             @������������������������       �                     �?0       1                    j�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK3KK&��hH�B�<        �?       @      �?      @      @      �?              �?                      �?                                      �?       @      �?       @              �?       @      �?                      �?      �?              �?       @              �?      �?      �?      �?      @      �?       @      �?       @      �?      @      @      �?              �?                      �?                                      �?       @      �?       @              �?       @      �?                      �?      �?              �?       @              �?      �?      �?      �?              �?       @      �?       @      �?      @                              �?                                                                                                                                                                      �?                                                                              �?              �?      @                              �?                                                                                                                                                                      �?                                                                              �?              �?                                      �?                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                              �?                                                                              �?              �?                                      �?                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                              �?                                      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                      @      �?                                      �?                                      �?       @      �?       @              �?       @      �?                      �?      �?                       @              �?      �?      �?      �?              �?       @                                      @      �?                                      �?                                                      �?       @                              �?                              �?                                                                                                                                      �?                                      �?                                                      �?       @                              �?                              �?                                                                                                                                      �?                                      �?                                                      �?                                      �?                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                      �?                                                                                              �?                                      �?                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                      �?                                                                                              �?                                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                      �?                                                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                                                                      �?       @                              �?       @                              �?                               @              �?      �?      �?      �?              �?       @                                                                                                                                                                               @                              �?                               @              �?                                                                                                                                                                                                                                                              �?                               @              �?                                                                                                                                                                                                                                                              �?                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                              �?       @                              �?                                                                                              �?      �?      �?              �?       @                                                                                                                              �?       @                              �?                                                                                                                                                                                                                                                                      �?                                      �?                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                                                                                              �?      �?      �?              �?       @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                      �?      �?      �?              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?      �?      �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                      �?              �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                      @                �t�bub��     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJ$�phG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hKhcK-hdh*h-K ��h/��R�(KK-��hk�B�	         ,                    l�@�A+K&:�?             C@       +                    f�@h+�v:�?             A@                           ̞@�&�'+�?             ?@������������������������       �                      @                            B�@��\P8�?             =@                           �@�?�'�@�?             3@                           �@������?             @       	                    ֞@      �?             @������������������������       �                     �?
                           ޞ@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           ��@      �?	             (@������������������������       �                      @                           �@��Q���?             $@                           
�@      �?             @                            �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �@9��8���?             @������������������������       �                      @                            �@      �?             @������������������������       �                     �?                           (�@VUUUUU�?             @������������������������       �                     �?                           4�@      �?              @������������������������       �                     �?������������������������       �                     �?!       "                    J�@�������?             $@������������������������       �                     @#       $                    N�@4և����?             @������������������������       �                      @%       (                    ^�@
ףp=
�?             @&       '                    V�@�q�q�?             @������������������������       �                     �?������������������������       �                      @)       *                    b�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK-KK&��hH�Bp5                �?      �?      �?       @              �?                      �?               @              �?      �?      �?       @      �?              �?      @                                              @               @      �?       @              @      �?              @      �?       @              �?      �?      �?       @              �?                      �?               @              �?      �?      �?       @      �?              �?      @                                              @               @      �?       @              @      �?                      �?       @              �?      �?      �?       @              �?                      �?               @              �?      �?      �?       @      �?              �?      @                                              @               @      �?       @                      �?                      �?       @                                                                                                                                                                                                                                       @                                                                                      �?      �?      �?       @              �?                      �?               @              �?      �?      �?       @      �?              �?      @                                              @                      �?       @                      �?                      �?       @              �?      �?      �?       @              �?                      �?               @              �?      �?      �?              �?                                                                      @                      �?       @                                                                      �?      �?      �?                                              �?                                                                                                                                      @                                                                                                      �?      �?      �?                                              �?                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                      �?              �?                                              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                              �?                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                                                                      @                                                                                                                               @              �?                                       @              �?      �?      �?              �?                                                                                              �?       @                                                                                                                                                       @                                                                                                                                                                                                                                                       @              �?                                                      �?      �?      �?              �?                                                                                              �?       @                                                                                               @              �?                                                                                      �?                                                                                                                                                                                                                      �?                                                                                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                                      �?      �?      �?                                                                                                              �?       @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                      �?      �?      �?                                                                                                              �?                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                      �?              �?                                                                                                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                              �?                                                                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                       @                      �?      @                                                                                                      �?                      �?       @                                                                                                                                                                      @                                                                                                                                                                                                                                                                               @                      �?                                                                                                              �?                      �?       @                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                      �?                                                                                                              �?                      �?       @                                                                                                                                                              �?                                                                                                                                               @                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                              �?                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                      @                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJW:+LhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hK
hcK-hdh*h-K ��h/��R�(KK-��hk�B�	                             
�@f��.�?             C@                           �@^N��)x�?             ,@                           ��@0�����?             "@       	                    �@4և����?             @                           �@      �?             @                           ؞@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @
                           ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                           �@�������?             8@������������������������       �                      @       ,                    n�@�����|�?             6@       +                    j�@H�z�G�?             4@       *                    f�@��^B{	�?             2@       !                    :�@     ��?             0@                           �@~X�<��?             "@                           �@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           &�@9��8���?             @                           �@VUUUUU�?             @������������������������       �                     �?                           "�@      �?              @������������������������       �                     �?������������������������       �                     �?                            *�@�q�q�?             @������������������������       �                      @������������������������       �                     �?"       #                    L�@������?             @������������������������       �                     @$       %                    R�@      �?             @������������������������       �                     �?&       '                    Z�@VUUUUU�?             @������������������������       �                     �?(       )                    b�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @�t�bh�h*h-K ��h/��R�(KK-KK&��hH�Bp5                                �?      �?      @              �?                               @       @      �?                               @       @      �?      @              �?                       @       @      �?              �?      �?      �?       @      �?       @       @      �?                                      �?              @              �?                               @                                               @                                      �?                               @                                                                                                                      �?                              �?                               @                                               @                                      �?                               @                                                                                                                      �?                              �?                               @                                                                                      �?                               @                                                                                                                      �?                              �?                                                                                                                                                       @                                                                                                                      �?                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                       @                                                                                      �?                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                      �?                                                               @      �?                                       @      �?      @                                       @              �?              �?      �?      �?       @      �?       @       @      �?                                                                                                                                                               @                                                                                                                                                                                              �?                                                               @      �?                                              �?      @                                       @              �?              �?      �?      �?       @      �?       @       @      �?                                              �?                                                               @      �?                                              �?      @                                       @              �?              �?      �?      �?       @      �?       @              �?                                              �?                                                               @      �?                                              �?      @                                       @              �?              �?      �?      �?       @      �?                      �?                                              �?                                                               @      �?                                              �?      @                                       @              �?              �?      �?      �?              �?                      �?                                              �?                                                               @      �?                                                                                               @                              �?      �?      �?                                                                                      �?                                                               @                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                      �?                                                                                               @                              �?      �?      �?                                                                                                                                                              �?                                                                                                                                      �?      �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                      �?                                                                                                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                               @                              �?                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                              �?      @                                                      �?                                              �?                      �?                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                      �?                                                              �?                                              �?                      �?                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                              �?                                              �?                      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                              �?                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                       @                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJF<KdhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hKhcK-hdh*h-K ��h/��R�(KK-��hk�B�	         $                    L�@�5��P�?             C@                           *�@!��w���?             =@                           "�@H�z�G�?             4@                           Ξ@�6�i�?             .@������������������������       �                      @                           �@�B�����?             *@                           
�@)\���(�?	             $@       	                    ڞ@      �?              @������������������������       �                     �?
                           �@ܶm۶m�?             @������������������������       �                     �?                           �@�������?             @������������������������       �                     �?                           �@�������?             @������������������������       �                     �?                           ��@      �?             @������������������������       �                     �?                           �@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           &�@���Q��?             @������������������������       �                     @������������������������       �                      @                           4�@��"e���?             "@������������������������       �                     @        !                    @�@�8��8��?             @������������������������       �                     @"       #                    F�@�q�q�?             @������������������������       �                     �?������������������������       �                      @%       &                    R�@�2�tk~�?             "@������������������������       �                     @'       (                    \�@�q�q�?             @������������������������       �                      @)       *                    h�@      �?             @������������������������       �                      @+       ,                    n�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK-KK&��hH�Bp5                �?                              �?      �?      �?      �?      �?      �?               @      @              @                       @      @       @                              �?       @      �?       @       @      @              �?               @      �?      �?                              �?                              �?      �?      �?      �?      �?      �?               @      @              @                       @               @                              �?       @      �?               @      @              �?                                                              �?                              �?      �?      �?      �?      �?      �?               @      @                                       @                                                       @      �?               @                      �?                                                              �?                              �?      �?      �?      �?      �?      �?               @                                               @                                                              �?               @                      �?                                                                                                                                                                                                                                                                                       @                                                                                      �?                              �?      �?      �?      �?      �?      �?               @                                               @                                                              �?                                      �?                                                              �?                              �?      �?      �?      �?      �?      �?                                                               @                                                              �?                                                                                                      �?                              �?      �?      �?      �?      �?      �?                                                                                                                              �?                                                                                                                                                      �?                                                                                                                                                                                                                                                              �?                              �?      �?              �?      �?      �?                                                                                                                              �?                                                                                                      �?                                                                                                                                                                                                                                                                                                                                              �?      �?              �?      �?      �?                                                                                                                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                      �?      �?              �?      �?                                                                                                                                      �?                                                                                                                                                                      �?                                                                                                                                                                                                                                                                              �?      �?              �?                                                                                                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                      �?      �?              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                      �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                               @                                                                                                                                                      �?                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                              @                                                                                               @                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                              @                                       @                              �?                                      @                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                              @                                       @                              �?                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                                                       @                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                      @                                                               @                                               @      �?      �?                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                                               @                                               @      �?      �?                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                               @      �?      �?                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                      �?      �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                      �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJؽ�hG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hK
hcK5hdh*h-K ��h/��R�(KK5��hk�B�                             Ξ@��D��?             C@                           ʞ@      �?             @������������������������       �                     �?������������������������       �                     @                           �@DSbq���?             A@                           ��@�z�G��?             $@                           �@      �?              @                           �@9��8���?             @	       
                    ֞@      �?             @������������������������       �                     �?                           ޞ@VUUUUU�?             @������������������������       �                     �?                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @                           �@      �?             8@                           �@4և����?             @                           �@
ףp=
�?             @                           
�@      �?              @������������������������       �                     �?������������������������       �                     �?                           �@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @                            $�@ҳ�wY;�?             1@                           �@�q�q�?             @������������������������       �                     �?������������������������       �                      @!       *                    N�@/�����?             ,@"       )                    H�@4և����?             @#       (                    >�@
ףp=
�?             @$       %                    *�@VUUUUU�?             @������������������������       �                     �?&       '                    2�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @+       ,                    R�@����X�?             @������������������������       �                      @-       .                    Z�@�������?             @������������������������       �                     �?/       0                    b�@      �?             @������������������������       �                     �?1       2                    f�@VUUUUU�?             @������������������������       �                     �?3       4                    l�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK5KK&��hH�B�>        @      �?      �?      �?       @      �?                               @      �?              �?              �?               @       @      �?       @              �?                       @      �?       @      �?      �?      �?       @       @      �?      �?              �?      �?              @                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                              @                                                                                                                                                                                                                                                                                                                      �?      �?      �?       @      �?                               @      �?              �?              �?               @       @      �?       @              �?                       @      �?       @      �?              �?       @       @      �?      �?              �?      �?                      �?      �?      �?                                               @      �?                                                       @                                                                       @                                                                                                      �?      �?      �?                                               @      �?                                                                                                                               @                                                                                                      �?      �?      �?                                               @      �?                                                                                                                                                                                                                                      �?      �?      �?                                                      �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?              �?                                                      �?                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                              �?                                                                      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                       @                                                                                                                                                                                                       @      �?                                                      �?              �?               @              �?       @              �?                       @      �?              �?              �?       @       @      �?      �?              �?      �?                                               @      �?                                                      �?                                              �?                                                                                               @                                                                                               @      �?                                                      �?                                              �?                                                                                                                                                                                                      �?                                                                                                      �?                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                               @                                                              �?                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                              �?               @                       @              �?                       @      �?              �?              �?               @      �?      �?              �?      �?                                                                                                                              �?                                                                                                                                       @                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                       @                       @              �?                       @      �?              �?              �?                      �?      �?              �?      �?                                                                                                                                               @                                      �?                       @      �?                              �?                                                                                                                                                                                                                                              �?                       @      �?                              �?                                                                                                                                                                                                                                              �?                              �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                       @                                                              �?                                      �?      �?              �?      �?                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                                                                                              �?                                      �?      �?              �?      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                      �?      �?              �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?      �?              �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                      �?                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                      �?                �t�bub��     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJX��vhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hKhcK5hdh*h-K ��h/��R�(KK5��hk�B�         2                    j�@�|�ʒ��?             C@                           ��@�E��'s�?             A@       
                    �@      �?              @                           ֞@
ףp=
�?             @                           Ξ@�q�q�?             @������������������������       �                     �?������������������������       �                      @       	                    ޞ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �@	j*D�?             :@                           �@�Q����?             @                           ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �@y'�L��?             5@                           �@�q�q�?             @                           �@      �?             @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           (�@�*;L�?             .@                           "�@�q�q�?             @������������������������       �                     �?������������������������       �                      @       #                    :�@9��8���?             (@       "                    4�@      �?             @        !                    .�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @$       %                    @�@      �?              @������������������������       �                     �?&       '                    F�@ܶm۶m�?             @������������������������       �                     �?(       )                    L�@�������?             @������������������������       �                     �?*       +                    V�@�������?             @������������������������       �                     �?,       -                    ^�@      �?             @������������������������       �                     �?.       /                    b�@VUUUUU�?             @������������������������       �                     �?0       1                    f�@      �?              @������������������������       �                     �?������������������������       �                     �?3       4                    n�@      �?             @������������������������       �                     @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK5KK&��hH�B�>        �?      �?       @      �?      �?                              �?                              �?       @       @      �?              �?      @      �?      �?       @              �?      �?              @                      �?       @      �?      �?      �?      @      �?      �?      �?      �?      �?       @      �?      �?                              �?                              �?       @       @      �?              �?      @      �?      �?       @              �?      �?              @                      �?       @      �?      �?      �?                      �?      �?      �?      �?       @      �?                                                                                                                                                                                      @                                                                                              �?      �?       @      �?                                                                                                                                                                                                                                                                                      �?               @                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                      �?              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      @                                                                                                                              �?                              �?                              �?       @       @      �?              �?      @      �?      �?       @              �?      �?                                      �?       @      �?      �?      �?                      �?      �?                                                                      �?                                                                      �?      @                                                                                                                                                                                                                              �?                                                                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                              �?                                                              �?       @       @      �?                              �?      �?       @              �?      �?                                      �?       @      �?      �?      �?                      �?      �?                                      �?                                                              �?               @                                                                                                                               @                                                                                              �?                                                              �?                                                                                                                                               @                                                                                              �?                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                       @              �?                              �?      �?       @              �?      �?                                      �?              �?      �?      �?                      �?      �?                                                                                                               @                                                                                                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                              �?                              �?      �?       @              �?      �?                                      �?                      �?      �?                      �?      �?                                                                                                                                                                               @              �?                                              �?                                                                                                                                                                                                                                                              �?                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                              �?                              �?      �?                              �?                                                              �?      �?                      �?      �?                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                              �?      �?                              �?                                                              �?      �?                      �?      �?                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                      �?      �?                                                                                              �?      �?                      �?      �?                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                      �?                                                                                                      �?      �?                      �?      �?                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                                      �?      �?                      �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                      �?      �?                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                              @      �?                                                                                                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                      �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���EhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hKhcK3hdh*h-K ��h/��R�(KK3��hk�B(                              �@��Ł�r�?             C@                           �@����%�?             3@                           ܞ@/�����?             ,@                           О@�q�q�?             @������������������������       �                     �?������������������������       �                      @       
                    �@N�zv�?	             &@       	                    �@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �@      �?              @                           �@      �?             @������������������������       �                     �?                           ��@VUUUUU�?             @������������������������       �                     �?                            �@      �?              @������������������������       �                     �?������������������������       �                     �?                           �@      �?             @������������������������       �                      @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?                           �@���Q��?             @������������������������       �                     @������������������������       �                      @                           &�@5mvq`��?             3@������������������������       �                     @                           2�@�6�i�?             .@������������������������       �                      @       &                    N�@�B�����?             *@        %                    J�@
ףp=
�?             @!       "                    @�@VUUUUU�?             @������������������������       �                     �?#       $                    F�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @'       ,                    ^�@      �?              @(       +                    X�@      �?             @)       *                    R�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @-       .                    b�@      �?             @������������������������       �                     �?/       0                    h�@VUUUUU�?             @������������������������       �                     �?1       2                    n�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK3KK&��hH�B�<        �?                              �?       @      �?       @               @      �?      �?      �?      @       @      �?       @      �?              �?      �?                              �?       @      �?      �?                      @                      �?      �?      �?      �?       @      �?                              �?       @      �?       @               @      �?      �?      �?               @                      �?                                                                      �?                              @                                                              �?                              �?       @      �?       @               @      �?      �?      �?                                      �?                                                                      �?                                                                                              �?                                                       @                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                      �?       @      �?                       @      �?      �?      �?                                      �?                                                                      �?                                                                                                                                                                       @      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                      �?       @      �?                                      �?      �?                                      �?                                                                      �?                                                                                                                                              �?                                      �?                                              �?                                                                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                              �?                                      �?                                              �?                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                      �?                                                                                      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                              �?       @                                                      �?                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                                      �?                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                               @                                                                                                                              @                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                      @              �?       @                      �?      �?                              �?       @              �?                                              �?      �?      �?      �?       @                                                                                                              @                                                                                                                                                                                                                                                                                                                              �?       @                      �?      �?                              �?       @              �?                                              �?      �?      �?      �?       @                                                                                                                                                                                                               @                                                                                                                                                                                                                              �?       @                      �?      �?                              �?                      �?                                              �?      �?      �?      �?       @                                                                                                                              �?       @                              �?                              �?                                                                                                                                                                                                                                      �?                                      �?                              �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                      �?                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                                                      �?                                                              �?                                              �?      �?      �?      �?       @                                                                                                                                                              �?                                                              �?                                                                               @                                                                                                                                                              �?                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                              �?      �?      �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                      �?      �?      �?                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                      �?      �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                      �?                �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ:9)bhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hK	hcK+hdh*h-K ��h/��R�(KK+��hk�Bh	         $                    R�@LM�]�?             C@                           �@�t�@��?             >@                           �@�.k���?
             1@                           �@�	j*D�?             *@                           ��@�z�G��?             $@                           ��@      �?              @       
                    �@9��8���?             @       	                    ڞ@      �?              @������������������������       �                     �?������������������������       �                     �?                           �@      �?             @������������������������       �                      @                           ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @                           �@      �?             @������������������������       �                     @������������������������       �                     �?                           �@ƵHPS!�?             *@������������������������       �                     @                           "�@0�����?             "@������������������������       �                     @                           ,�@�������?             @������������������������       �                     �?                           6�@�������?             @������������������������       �                     �?                           @�@      �?             @������������������������       �                     �?        !                    F�@VUUUUU�?             @������������������������       �                     �?"       #                    L�@      �?              @������������������������       �                     �?������������������������       �                     �?%       &                    X�@      �?              @������������������������       �                     @'       (                    ^�@�Q����?             @������������������������       �                     @)       *                    d�@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK+KK&��hH�B3                        �?                              @               @              �?      �?      �?              @      �?               @      @      �?      �?              �?      �?      �?      �?       @      @                      @              �?                              �?      @                      �?                              @               @              �?      �?      �?              @      �?               @      @      �?      �?              �?      �?      �?      �?       @                              @                                                                              �?                              @               @              �?      �?      �?                                       @      @                              �?                               @                                                                                                              �?                              @               @              �?      �?                                               @                                      �?                               @                                                                                                              �?                                               @              �?      �?                                               @                                      �?                               @                                                                                                              �?                                                              �?      �?                                               @                                      �?                               @                                                                                                              �?                                                              �?      �?                                                                                      �?                               @                                                                                                              �?                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                      �?                                                                                      �?                               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                      �?                                                                                      �?                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                              �?                                              @                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                              @      �?                              �?      �?                      �?      �?      �?                                      @                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                              @      �?                              �?      �?                      �?      �?      �?                                                                                                                                                                                                                      @                                                                                                                                                                                                                                                                                                                      �?                              �?      �?                      �?      �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                              �?                              �?      �?                      �?      �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                              �?                              �?      �?                              �?                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                              �?      �?                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                      �?      �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                      �?                                                                                                                                                                                                                                                                                                                                                                              @                                      �?                              �?      @                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                      �?                              �?      @                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                      �?                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                              �?                                        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�BHzhG        hNhG        h%Kh&Kh'h*h-K ��h/��R�(KK&��hH�B0                �?       @      @      @      @      @      @       @      "@      $@      &@      (@      *@      ,@      .@      0@      1@      2@      3@      4@      5@      6@      7@      8@      9@      :@      ;@      <@      =@      >@      ?@      @@     �@@      A@     �A@      B@     �B@�t�bh<hMhPC&       ���R�hUKhVhYKh*h-K ��h/��R�(KK��hP�C&       �t�bK��R�}�(hKhcK)hdh*h-K ��h/��R�(KK)��hk�B�                             ֞@�� 'a��?             C@������������������������       �                     @       (                    f�@      �?             @@                           ��@��\P8�?             =@       
                    ��@����>4�?             @                           ޞ@      �?             @������������������������       �                      @       	                    �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �@���|���?             6@������������������������       �                      @       '                    `�@q=
ףp�?             4@       &                    X�@l~X�<�?             2@                            �@      �?             0@                           �@�q�q�?             @                           �@      �?             @                           �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @       !                    >�@��Q���?             $@                           .�@9��8���?             @                           &�@VUUUUU�?             @������������������������       �                     �?                           *�@      �?              @������������������������       �                     �?������������������������       �                     �?                            4�@�q�q�?             @������������������������       �                      @������������������������       �                     �?"       #                    J�@      �?             @������������������������       �                      @$       %                    R�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK)KK&��hH�B�0                �?      @       @      �?                               @                      �?              �?       @                              �?      �?              �?      @       @       @      �?              �?              �?       @              @       @                               @                      @                                                                                                                                                                                                                                                                                                      �?               @      �?                               @                      �?              �?       @                              �?      �?              �?      @       @       @      �?              �?              �?       @              @       @                               @              �?               @      �?                               @                      �?              �?       @                              �?      �?              �?      @       @       @      �?              �?              �?       @                       @                               @              �?               @                                                              �?                                                                                      @                                                                                                                                      �?               @                                                              �?                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                              �?                                                                              �?                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                      @                                                                                                                                                              �?                               @                                      �?       @                              �?      �?              �?               @       @      �?              �?              �?       @                       @                               @                                                                       @                                                                                                                                                                                                                                                                              �?                                                                      �?       @                              �?      �?              �?               @       @      �?              �?              �?       @                       @                               @                                      �?                                                                      �?       @                              �?      �?              �?               @       @      �?              �?              �?       @                                                       @                                      �?                                                                      �?       @                              �?      �?              �?               @       @      �?              �?              �?       @                                                                                              �?                                                                               @                              �?                                                                                               @                                                                                              �?                                                                                                              �?                                                                                               @                                                                                              �?                                                                                                              �?                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                      �?                                              �?              �?               @       @      �?              �?              �?                                                                                                                                                                              �?                                                              �?               @              �?                              �?                                                                                                                                                                              �?                                                                                              �?                              �?                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                                              �?                              �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                              �?               @                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                              �?                                       @                      �?                                                                                                                                                                                                                                                                                       @                                                                                                                                                                                                                                                                      �?                                                              �?                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                              �?                                                                                                                                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                               @                                                                                                                                                                                                                                                                                                      @                                        �t�bub�       hhubehhub.